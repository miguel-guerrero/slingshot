//----------------------------------------------------------------------------
// adder
//----------------------------------------------------------------------------
module adder 
#(
    parameter W = 8)
(
    input [7999:0] ins,
    output reg [W+1:0] sm
);




always @(*) begin : combo_logic
    sm = ins/*[1,1][9,4,1]*/[7999:7980];
end


endmodule


