//----------------------------------------------------------------------------
// adder
//----------------------------------------------------------------------------
module adder 
#(
    parameter W = 8)
(
    input [1999:0] ins,
    output reg [W+1:0] sm
);




always @(*) begin : combo_logic
    sm = ins/*[9,4,1]*/[1999:1980];
end


endmodule


